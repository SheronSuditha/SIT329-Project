module volts_to_temp (
	input voltage
);

endmodule